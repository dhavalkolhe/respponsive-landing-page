/mnt/c/users/dhava/Desktop/Web-dev/responsove-headphone-landing-page